`ifndef GLOBAL_PARAMS_VH
`define GLOBAL_PARAMS_VH


`define  ADD 4'b0010;
`define  SUB 4'b0110;
`define  AND 4'b0000;
`define  OR  4'b0001;
`define  XOR 4'b0100;
`define  SLL 4'b0101; // Shift left logical
`define  SRL 4'b0110; // Shift right logical
`define  SRA 4'b0111; // Shift right arithmetic


`endif